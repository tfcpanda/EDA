module MUX41a2 (A, B, C, D, S1, S0, Y);